module Bus(bus);
    input wand bus;

    assign bus = 'b1;
    
endmodule