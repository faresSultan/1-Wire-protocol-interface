module Bus(bus);
    inout wand bus;

    assign bus = 'b1;
    
endmodule